
// This file contains multiple modules. 
//   Verilator likes 1 file for each module
/* verilator lint_off DECLFILENAME */
/* verilator lint_off UNUSED */
/* verilator lint_off BLKSEQ */
/* verilator lint_off WIDTH */

// Include Vmicro16 ISA containing definitions for the bits
`include "vmicro16_isa.v"

// This module aims to be a SYNCHRONOUS, WRITE_FIRST BLOCK RAM
//   https://www.xilinx.com/support/documentation/user_guides/ug473_7Series_Memory_Resources.pdf
//   https://www.xilinx.com/support/documentation/user_guides/ug383.pdf
//   https://www.xilinx.com/support/documentation/sw_manuals/xilinx2016_4/ug901-vivado-synthesis.pdf
module vmicro16_bram # (
        parameter MEM_WIDTH    = 16,
        parameter MEM_DEPTH    = 256
) (
        input clk, input reset,
        
        input      [MEM_WIDTH-1:0] mem_addr,
        input      [MEM_WIDTH-1:0] mem_in,
        input                      mem_we,
        output reg [MEM_WIDTH-1:0] mem_out
);
        // memory vector
        reg [MEM_WIDTH-1:0] mem [0:MEM_DEPTH-1];

        // not synthesizable
        integer i;
        initial for (i = 0; i < MEM_DEPTH; i = i + 1) mem[i] <= 0;

        always @(posedge clk) begin
                // synchronous WRITE_FIRST (page 13)
                if (mem_we) begin
                        mem[mem_addr] <= mem_in;
                        $display($time, "\tbram: W mem[%h] <= %h", mem_addr, mem_in);
                end else begin
                        mem_out <= mem[mem_addr];
                end
        end

        // TODO: Reset impl = every clock while reset is asserted, clear each cell
        //       one at a time, mem[i++] <= 0
endmodule

// Wishbone wrapper around the register file to use as a peripheral
module vmicro16_regs_wb # (
        parameter CELL_WIDTH    = 16,
        parameter CELL_DEPTH    = 8,
        parameter CELL_SEL_BITS = 3,
        parameter CELL_DEFAULTS = 0,
        parameter DEBUG_NAME    = "",
        parameter PIPELINE_READ = 0
) (
        input clk, input reset,

        // wishbone slave interface
        input                   wb_stb_i,
        input                   wb_cyc_i,
        input                   wb_we_i,
        input  [CELL_WIDTH-1:0] wb_addr_i,
        input  [CELL_WIDTH-1:0] wb_data_i,
        output [CELL_WIDTH-1:0] wb_data_o,
        output                  wb_ack_o,
        output                  wb_stall_o,
        output                  wb_err_o
);
        // embedded register data
        wire [CELL_SEL_BITS-1:0] reg_rs1;
        wire [CELL_WIDTH-1:0]    reg_rd1;
        wire                     reg_we;
        wire [CELL_WIDTH-1:0]    reg_wd;

        reg selected;
        always @(*) begin
                if (wb_stb_i) 
                        selected = 1'b1;
                else if (selected && wb_cyc_i)
                        selected = 1'b1;
                else if (selected && !wb_cyc_i) 
                        selected = 1'b0;
                else    selected = 1'b0;
        end

        assign reg_we  = wb_we_i && wb_stb_i;
        assign reg_rs1 = wb_addr_i[CELL_SEL_BITS-1:0];
        assign reg_wd  = wb_data_i;
        
        // Only stall on write requests
        //assign wb_stall_o = wb_cyc_i && wb_we_i;
        // TODO: Stall for 1 clock if pipelined
        assign wb_stall_o = PIPELINE_READ ? wb_stb_i : 1'b0;
        // Only use the output bus when we're selected and it's a read req
        assign wb_data_o  = (selected && !wb_we_i)    ? reg_rd1 : {(CELL_WIDTH-1){1'bZ}};
        // TODO: ack on same stb clock allowed?
        assign wb_ack_o   = (wb_cyc_i && !wb_stall_o) ? 1'b1 : 1'bZ;

        vmicro16_regs # (
                .CELL_WIDTH     (CELL_WIDTH),
                .CELL_DEPTH     (CELL_DEPTH),
                .CELL_SEL_BITS  (CELL_SEL_BITS),
                .CELL_DEFAULTS  (CELL_DEFAULTS),
                .DEBUG_NAME     (DEBUG_NAME),
                .PIPELINE_READ  (PIPELINE_READ)
        ) vmicro16_regs_wb_i (
                 .clk           (clk)
                ,.reset         (reset)
                // Read port 1 (IDEX)
                ,.rs1           (reg_rs1)
                ,.rd1           (reg_rd1)
                // Read port 2 (IDEX) unused
                //,.rs2           (dec_rs2)
                //,.rd2           (reg_rd2)
                // Write port (MEWB)
                ,.we            (reg_we)
                ,.ws1           (reg_rs1)
                ,.wd            (reg_wd)
        );
endmodule

module vmicro16_regs # (
        parameter CELL_WIDTH    = 16,
        parameter CELL_DEPTH    = 8,
        parameter CELL_SEL_BITS = 3,
        parameter CELL_DEFAULTS = 0,
        parameter DEBUG_NAME    = "",
        parameter PIPELINE_READ = 0
) (
        input clk, input reset,
        // ID/EX stage reg reads
        // Dual port register reads
        input      [CELL_SEL_BITS-1:0] rs1, // port 1
        output reg [CELL_WIDTH-1:0]    rd1,
        input      [CELL_SEL_BITS-1:0] rs2, // port 2
        output reg [CELL_WIDTH-1:0]    rd2,
        // EX/WB final stage write back
        input                          we,
        input [CELL_SEL_BITS-1:0]      ws1,
        input [CELL_WIDTH-1:0]         wd
);
        reg [CELL_WIDTH-1:0] regs [0:CELL_DEPTH-1] /*verilator public_flat*/;
        
        // Initialise registers with default values
        //   Really only used for special registers used by the soc
        // TODO: How to do this on reset?
        initial if (CELL_DEFAULTS) $readmemh(CELL_DEFAULTS, regs);

        integer i;
        always @(posedge clk) 
                if (reset) 
                        if (CELL_DEFAULTS) $readmemh(CELL_DEFAULTS, regs); // TODO:
                        else for(i = 0; i < CELL_DEPTH; i = i + 1) regs[i] <= {(CELL_WIDTH-1){1'b0}}; 
                else if (we) begin
                        $display($time, "\tREGS #%s: Writing %h to reg[%d]", DEBUG_NAME, wd, ws1);
                        $display($time, "\t\t\t| %h %h %h %h | %h %h %h %h |", 
                                regs[0], regs[1], regs[2], regs[3], regs[4], regs[5], regs[6], regs[7]);
                        // Perform the right
                        regs[ws1] <= wd;
                end

        generate if (PIPELINE_READ) 
                always @(posedge clk) 
                        if (reset) begin
                                rd1 <= {(CELL_WIDTH-1){1'b0}};
                                rd2 <= {(CELL_WIDTH-1){1'b0}};
                        end else begin
                                rd1 <= regs[rs1];
                                rd2 <= regs[rs2];
                        end
        else
                always @(*) begin
                        rd1 = regs[rs1];
                        rd2 = regs[rs2];
                end
        endgenerate
endmodule

// Decoder is hard to parameterise as it's very closely linked to the ISA.
module vmicro16_dec # (
        parameter INSTR_WIDTH    = 16,
        parameter INSTR_OP_WIDTH = 5,
        parameter INSTR_RS_WIDTH = 3,
        parameter ALU_OP_WIDTH   = 5
) (
        //input clk,   // not used yet (all combinational)
        //input reset, // not used yet (all combinational)

        input  [INSTR_WIDTH-1:0]    instr,

        output [INSTR_OP_WIDTH-1:0] opcode,
        output [INSTR_RS_WIDTH-1:0] rd,
        output [INSTR_RS_WIDTH-1:0] ra,
        output [7:0]                imm8,
        output [11:0]               imm12,
        output [4:0]                simm5,

        // This can be freely increased without affecting the isa
        output reg [ALU_OP_WIDTH-1:0] alu_op,

        output reg has_imm8,
        output reg has_imm12,
        output reg has_we,
        output reg has_br,
        output reg has_mem,
        output reg has_mem_we,

        output halt
        
        // TODO: Use to identify bad instruction and
        //       raise exceptions
        //,output     is_bad 
);
        assign opcode = instr[15:11];
        assign rd     = instr[10:8];
        assign ra     = instr[7:5];
        assign imm8   = instr[7:0];
        assign imm12  = instr[11:0];
        assign simm5  = instr[4:0];
        // Special opcodes
        assign halt   = (opcode == `VMICRO16_OP_HALT);

        // exme_op
        always @(*) case (opcode)
                `VMICRO16_OP_HALT, // TODO: stop ifid
                `VMICRO16_OP_NOP:             alu_op = `VMICRO16_ALU_NOP;
                
                `VMICRO16_OP_LW:              alu_op = `VMICRO16_ALU_LW;
                `VMICRO16_OP_SW:              alu_op = `VMICRO16_ALU_SW;

                `VMICRO16_OP_MOV:             alu_op = `VMICRO16_ALU_MOV;
                `VMICRO16_OP_MOVI:            alu_op = `VMICRO16_ALU_MOVI;
                `VMICRO16_OP_MOVI_L:          alu_op = `VMICRO16_ALU_MOVI_L; 

                `VMICRO16_OP_BR:              alu_op = `VMICRO16_ALU_BR;
                
                `VMICRO16_OP_BIT:         casez (simm5)
                        `VMICRO16_OP_BIT_OR:      alu_op = `VMICRO16_ALU_BIT_OR;
                        `VMICRO16_OP_BIT_XOR:     alu_op = `VMICRO16_ALU_BIT_XOR;
                        `VMICRO16_OP_BIT_AND:     alu_op = `VMICRO16_ALU_BIT_AND;
                        `VMICRO16_OP_BIT_NOT:     alu_op = `VMICRO16_ALU_BIT_NOT;
                        `VMICRO16_OP_BIT_LSHFT:   alu_op = `VMICRO16_ALU_BIT_LSHFT;
                        `VMICRO16_OP_BIT_RSHFT:   alu_op = `VMICRO16_ALU_BIT_RSHFT;
                        default:                  alu_op = `VMICRO16_ALU_BAD; endcase

                `VMICRO16_OP_ARITH_U:     casez (simm5)
                        `VMICRO16_OP_ARITH_UADD:  alu_op = `VMICRO16_ALU_ARITH_UADD;
                        `VMICRO16_OP_ARITH_USUB:  alu_op = `VMICRO16_ALU_ARITH_USUB;
                        `VMICRO16_OP_ARITH_UADDI: alu_op = `VMICRO16_ALU_ARITH_UADDI;
                        default:                  alu_op = `VMICRO16_ALU_BAD; endcase
                
                `VMICRO16_OP_ARITH_S:     casez (simm5)
                        `VMICRO16_OP_ARITH_SADD:  alu_op = `VMICRO16_ALU_ARITH_SADD;
                        `VMICRO16_OP_ARITH_SSUB:  alu_op = `VMICRO16_ALU_ARITH_SSUB;
                        `VMICRO16_OP_ARITH_SSUBI: alu_op = `VMICRO16_ALU_ARITH_SSUBI; 
                        default:                  alu_op = `VMICRO16_ALU_BAD; endcase
                
                default: begin
                        alu_op = `VMICRO16_ALU_BAD;
                        $display($time, "\tDEC: unknown opcode: %h", opcode);
                end
        endcase

        // Register writes
        always @(*) case (opcode)
                `VMICRO16_OP_LW,
                `VMICRO16_OP_MOV,
                `VMICRO16_OP_MOVI,
                `VMICRO16_OP_MOVI_L,
                `VMICRO16_OP_ARITH_U,
                `VMICRO16_OP_ARITH_S,
                `VMICRO16_OP_CMP,
                `VMICRO16_OP_SETC:          has_we = 1'b1;
                default:                    has_we = 1'b0;
        endcase

        // Contains 8-bit immediate
        always @(*) case (opcode)
                `VMICRO16_OP_MOVI,
                `VMICRO16_OP_CMP:           has_imm8 = 1'b1;
                default:                    has_imm8 = 1'b0;
        endcase

        // Contains 12-bit immediate
        always @(*) case (opcode)
                `VMICRO16_OP_MOVI_L:        has_imm12 = 1'b1;
                default:                    has_imm12 = 1'b0;
        endcase
        
        // Will branch the pc
        always @(*) case (opcode)
                `VMICRO16_OP_BR:            has_br = 1'b1;
                default:                    has_br = 1'b0;
        endcase
        
        // Requires external memory
        always @(*) case (opcode)
                `VMICRO16_OP_LW,
                `VMICRO16_OP_SW:            has_mem = 1'b1;
                default:                    has_mem = 1'b0;
        endcase
        
        // Requires external memory write
        always @(*) case (opcode)
                `VMICRO16_OP_SW:            has_mem_we = 1'b1;
                default:                    has_mem_we = 1'b0;
        endcase
endmodule


module vmicro16_alu # (
    parameter OP_WIDTH   = 5,
    parameter DATA_WIDTH = 16
) (
        // input clk, // TODO: make clocked

        input      [OP_WIDTH-1:0]   op,
        input      [DATA_WIDTH-1:0] d1, // rs1/dst
        input      [DATA_WIDTH-1:0] d2, // rs2
        output reg [DATA_WIDTH-1:0] q
);
        always @(*) case (op)
                `VMICRO16_ALU_BR,
                `VMICRO16_ALU_NOP:          q = 0;

                `VMICRO16_ALU_LW,
                `VMICRO16_ALU_SW:           q = d2;

                `VMICRO16_ALU_BIT_OR:       q = d1 | d2;
                `VMICRO16_ALU_BIT_XOR:      q = d1 ^ d2;
                `VMICRO16_ALU_BIT_AND:      q = d1 & d2;
                `VMICRO16_ALU_BIT_NOT:      q = ~(d2);
                `VMICRO16_ALU_BIT_LSHFT:    q = d1 << d2;
                `VMICRO16_ALU_BIT_RSHFT:    q = d1 >> d2;

                `VMICRO16_ALU_MOV:          q = d2;
                `VMICRO16_ALU_MOVI:         q = d2;
                `VMICRO16_ALU_MOVI_L:       q = d2;

                `VMICRO16_ALU_ARITH_UADD:   q = d1 + d2;
                `VMICRO16_ALU_ARITH_USUB:   q = d1 - d2;
                // TODO: ALU should have simm5 as input
                `VMICRO16_ALU_ARITH_UADDI:  q = d1 + d2;
                
                `VMICRO16_ALU_ARITH_SADD:   q = $signed(d1) + $signed(d2);
                `VMICRO16_ALU_ARITH_SSUB:   q = $signed(d1) - $signed(d2);
                // TODO: ALU should have simm5 as input
                `VMICRO16_ALU_ARITH_SSUBI:  q = $signed(d1) + $signed(d2);


                // TODO: Parameterise
                default: begin
                        $display($time, "\tALU: unknown op: %h", op);
                        q = {(DATA_WIDTH-1){1'bZZZZ}};
                end
        endcase
endmodule

module vmicro16_mewb (
        input clk,
        input reset,

        input [15:0] exme_pc,  output reg [15:0] mewb_pc,
        
        input [15:0] exme_d, 
        input [15:0] mem_out,  output reg [15:0] mewb_d,
        
        input [15:0] exme_d2,  output reg [15:0] mewb_d2,
        input [2:0]  exme_rs1, output reg [2:0]  mewb_rs1,

        input      [15:0] exme_jmp_target, 
        output reg [15:0] mewb_jmp_target,

        input exme_has_br,      output reg mewb_has_br,
        input exme_has_we,      output reg mewb_has_we,
        input exme_has_mem,     output reg mewb_has_mem,
        input exme_has_mem_we,  output reg mewb_has_mem_we,

        input valid_mem,
        input valid_stage1,     output reg valid_mewb,

        input jmping
);
        // MEWB stage
        always @(posedge clk)
        if (!reset) begin
                if (valid_stage1) begin
                        // Move previous stage regs into this stage
                        mewb_pc         <= exme_pc; // Only for simulation
                        
                        if (exme_has_mem) mewb_d <= mem_out;
                        else              mewb_d <= exme_d;
                        
                        mewb_d2         <= exme_d2;
                        mewb_rs1        <= exme_rs1;
                        mewb_jmp_target <= exme_jmp_target;

                        mewb_has_br      <= exme_has_br;
                        mewb_has_we      <= exme_has_we;
                        mewb_has_mem     <= exme_has_mem;
                        mewb_has_mem_we  <= exme_has_mem_we;
                        
                        if (exme_has_mem) 
                                if (exme_has_mem_we)
                                        $display($time, "\tmmu: SW: RAM[%h] <= r[%h] (%h)",
                                                exme_d, exme_rs1, exme_d2);
                                else
                                        $display($time, "\tmmu: LW: r[%h] <= RAM[%h]",
                                                exme_rs1, exme_d);
                end
                valid_mewb <= valid_stage1 && !jmping && valid_mem;
        end else begin
                valid_mewb      <= 1'b0;
                mewb_has_br     <= 1'b0;
                mewb_has_we     <= 1'b0;
                mewb_has_mem    <= 1'b0;
                mewb_has_mem_we <= 1'b0;
        end
endmodule

module vmicro16_wb (
        input clk,
        input reset,
        
        input jmping,

        input [15:0] mewb_d,          output reg [15:0] wb_d,
        input [2:0]  mewb_rs1,        output reg [2:0]  wb_rs1,
        input        mewb_has_we,     output reg        wb_we,
        input        mewb_has_br,     output reg        wb_has_br,
        input [15:0] mewb_jmp_target, output reg [15:0] wb_jmp_target,
        
        input valid_mewb,             output reg valid_wb
);
        // WB stage
        always @(posedge clk)
        if (!reset) begin
                if (valid_mewb) begin
                        wb_d          <= mewb_d;
                        wb_we         <= mewb_has_we;
                        wb_rs1        <= mewb_rs1;
                        wb_has_br     <= mewb_has_br;
                        wb_jmp_target <= mewb_jmp_target;
                end
                valid_wb <= valid_mewb && !jmping;
        end else begin
                valid_wb      <= 1'b0;
                wb_we         <= 1'b0;
                wb_has_br     <= 1'b0;
                wb_jmp_target <= 1'b0;
        end
endmodule


module vmicro16_mmu # (
        parameter MEM_WIDTH    = 16,
        parameter MEM_DEPTH    = 1024,

        parameter MEM_RVAL     = 16'h00CC
) (
        input clk,
        input reset,

        output valid,

        input req,

        input  [15:0] mem_addr,
        input  [15:0] mem_in,
        input         mem_we,
        input  [1:0]  mem_whl, // TODO: apply to mem_out
        output reg [15:0] mem_out,

        // wishbone peripheral master
        output reg    wb_mosi_stb_o_regs,
        //output wb_stb_o_xx,
        output reg    wb_mosi_cyc_o,
        output [15:0] wb_mosi_addr_o,
        output        wb_mosi_we_o,
        output [15:0] wb_mosi_data_o, // seperate data_o and data_i buses
        input  [15:0] wb_miso_data_i, // seperate data_o and data_i buses
        
        input         wb_miso_ack_i
);
        wire [15:0] bram_out;

        ////////////////////////////////
        //        TODO: CLEANUP
        ////////////////////////////////
        reg active = 0;
        always @(*)
        if (req) begin
                active = 1'b1;
        end else if (wb_miso_ack_i) begin
                active = 1'b0;
        end else 
                active = active;

        ////////////////////////////////
        //        TODO: CLEANUP
        ////////////////////////////////
        always @(*)
        if (reset) 
                mem_out = 16'h0;
        else if(active && wb_mosi_stb_o_regs) begin
                wb_mosi_cyc_o = 1'b1;
                if (wb_miso_ack_i) begin
                        mem_out = wb_miso_data_i;
                end
        end else if (active) begin
                mem_out = bram_out;
        end else begin
                wb_mosi_cyc_o = 1'b0;
                // TODO: mem_out isn't valid in this state, output high z or 0?
                mem_out = 16'hZZ;
        end

        // bram memory is always single clk, wb is unknown
        assign valid = active ? wb_miso_ack_i : 1'b1;

        ////////////////////////////////
        //        TODO: CLEANUP
        ////////////////////////////////
        // Virtual memory translator
        always @(*) begin
                // zero all peripherals
                wb_mosi_stb_o_regs = 0;

                if (req) begin
                        // enable peripherals when their address is selected
                        casez(mem_addr)
                                15'h01??: wb_mosi_stb_o_regs = 1'b1;
                                default:  wb_mosi_stb_o_regs = 1'b0;
                        endcase
                end
        end

        wire   wb_active      = wb_mosi_cyc_o; // deprecated
        wire   wb_stb         = wb_mosi_stb_o_regs;// || req;
        //assign wb_mosi_cyc_o  = wb_stb;
        assign wb_mosi_we_o   = wb_active ? mem_we   : 1'b0;
        assign wb_mosi_addr_o = wb_active ? mem_addr : 16'h00;
        assign wb_mosi_data_o = wb_active ? mem_in   : 16'h00;

        //assign mem_out        = wb_active ? wb_miso_data_i : bram_out;


        // TODO: Should this be inside the mmu or outside?
        wire bram_we = mem_we && !wb_active;
        vmicro16_bram # (
                .MEM_WIDTH(MEM_WIDTH), // TODO: mem 16b or 8b wide?
                .MEM_DEPTH(MEM_DEPTH)
        ) bram (
                .clk            (clk), 
                .reset          (reset), 
                // port 1
                .mem_addr       (mem_addr), 
                .mem_in         (mem_in), 
                .mem_we         (bram_we), 
                .mem_out        (bram_out)
        );

        // reset must be held long for atleast MEM_SIZE clocks
        // to fully erase the bram. 
        //   E.g. Xilinx bram 1024 cells = 1024 clocks = ~21us
        // TODO: implement with a dfa
endmodule


module vmicro16_stage1new (
        input clk,
        input reset,
        input stall,
        
        // debug
        output reg [15:0] stage1_pc,

        output reg valid_stage1,

        // sync decoder outputs
        output reg [15:0] stage_instrc,
        output reg [4:0] stage1_op,
        output reg [2:0] stage1_rs1c,
        output reg [2:0] stage1_rs2c,
        output reg       stage1_has_imm8,
        output reg       stage1_has_simm5,
        output reg       stage1_has_we,
        output reg       stage1_has_br,
        output reg       stage1_has_mem,
        output reg       stage1_has_mem_we,
        output reg       stage1_halt,

        // sync ALU outputs
        output reg [15:0] stage1_alu_d,
        output reg [15:0] stage1_alu_d2,
        
        // async outputs
        output     [2:0] stage1_rs1,
        output     [2:0] stage1_rs2,

        // async register reads
        input      [15:0] reg_rd1,
        input      [15:0] reg_rd2
);

        reg [15:0] pc;
        initial pc = 0;

        // Instruction memory
        reg [7:0] mem_cache [0:31];
        integer i;
        // Initialise instruction memory
        initial begin
                $display($time, "\tResetting mem");
                for(i = 0; i < 32; i = i + 1) mem_cache[i] = 8'h00;
                
                /*
                // MOV 1 R0
                mem_cache[0]  = {`VMICRO16_OP_MOVI,    3'h0}; mem_cache[1]  = { 8'h01 };
                // ADDI 1 R0
                mem_cache[2]  = {`VMICRO16_OP_ARITH_U, 3'h0}; mem_cache[3]  = {3'h7, 1'b0, 4'h1};
                //*/

                //*
                // register dependency
                mem_cache[0]  = {`VMICRO16_OP_MOVI,    3'h5}; mem_cache[1]  = { 8'h01 };
                mem_cache[2]  = {`VMICRO16_OP_ARITH_U, 3'h5}; mem_cache[3]  = {3'h7, 1'b0, 4'h2};
                //*/

                /*
                // Single cycle register writes
                // Should execute 1 clock each
                mem_cache[0]  = {`VMICRO16_OP_MOVI, 3'h0}; mem_cache[1]  = { 8'h00 };
                mem_cache[2]  = {`VMICRO16_OP_MOVI, 3'h1}; mem_cache[3]  = { 8'h01 };
                mem_cache[4]  = {`VMICRO16_OP_MOVI, 3'h2}; mem_cache[5]  = { 8'h02 };
                mem_cache[6]  = {`VMICRO16_OP_MOVI, 3'h3}; mem_cache[7]  = { 8'h03 };
                mem_cache[8]  = {`VMICRO16_OP_MOVI, 3'h4}; mem_cache[9]  = { 8'h04 };
                mem_cache[10] = {`VMICRO16_OP_MOVI, 3'h5}; mem_cache[11] = { 8'h05 };
                mem_cache[12] = {`VMICRO16_OP_MOVI, 3'h6}; mem_cache[13] = { 8'h06 };
                mem_cache[14] = {`VMICRO16_OP_MOVI, 3'h7}; mem_cache[15] = { 8'h07 };
                mem_cache[16] = {`VMICRO16_OP_HALT, 3'h0}; mem_cache[17] = { 8'h00 };
                //*/
                
                /*
                // while (1) add loop
                mem_cache[0]  = {`VMICRO16_OP_MOVI,    3'h0}; mem_cache[1]  = { 8'h00 };
                mem_cache[2]  = {`VMICRO16_OP_MOVI,    3'h1}; mem_cache[3]  = { -8'd02 };
                mem_cache[4]  = {`VMICRO16_OP_ARITH_U, 3'h0}; mem_cache[5]  = {3'h7, 1'b0, 4'h1};
                mem_cache[6]  = {`VMICRO16_OP_ARITH_U, 3'h0}; mem_cache[7]  = {3'h7, 1'b0, 4'h3};
                mem_cache[8]  = {`VMICRO16_OP_ARITH_U, 3'h0}; mem_cache[9]  = {3'h7, 1'b0, 4'h5};
                mem_cache[10] = {`VMICRO16_OP_BR,      3'h1}; mem_cache[11] = {`VMICRO16_OP_BR_U};
                mem_cache[12] = {`VMICRO16_OP_NOP,     3'h0}; mem_cache[13] = {8'h0};
                mem_cache[14] = {`VMICRO16_OP_NOP,     3'h0}; mem_cache[15] = {8'h0};
                mem_cache[16] = {`VMICRO16_OP_NOP,     3'h0}; mem_cache[17] = {8'h0};
                mem_cache[18] = {`VMICRO16_OP_NOP,     3'h0}; mem_cache[19] = {8'h0};
                mem_cache[20] = {`VMICRO16_OP_HALT,    3'h0}; mem_cache[21] = {8'h00};
                //*/
        end

        // Every clock:
        //   get new instruction
        //   decode instruction
        //   fetch operands
        //   alu it

        reg f_valid = 1;
        reg d_valid = 0;
        reg e_valid = 0;

        reg  [15:0] stage1_instr;
        always @(*) begin
                if (reset) begin
                        stage1_instr = 0;
                end else begin
                        // Load current instruction from memory
                        stage1_instr = {mem_cache[pc], mem_cache[pc+1]};
                end
        end

        always @(posedge clk) begin
                if (reset) begin
                        pc <= 0;
                        stage1_pc <= 0;

                        // Clock outputs
                        stage_instrc      <= 0;
                        stage1_pc         <= 0;
                        stage1_op         <= 0;
                        stage1_rs1c       <= 0;
                        stage1_rs2c       <= 0;
                        //stage1_imm8       <= 0;
                        stage1_has_imm8   <= 0;
                        //stage1_has_simm5  <= 0;
                        stage1_has_br     <= 0;
                        stage1_has_we     <= 0;
                        stage1_has_mem    <= 0;
                        stage1_has_mem_we <= 0;
                        //stage1_alu_op     <= 0;
                        stage1_halt       <= 0;
                        valid_stage1       <= 0;
                end
                else begin
                        if (!stall) begin
                                // Move to next instruction
                                pc        <= pc + 2;

                                // Clock outputs
                                stage_instrc      <= stage1_instr;
                                stage1_pc         <= pc;
                                stage1_op         <= w_stage1_op;
                                stage1_rs1c       <= stage1_rs1;
                                stage1_rs2c       <= stage1_rs2;
                                //stage1_imm8       <= w_stage1_imm8;
                                stage1_has_imm8   <= w_stage1_has_imm8;
                                //stage1_has_simm5  <= w_stage1_has_simm5;
                                stage1_has_br     <= w_stage1_has_br;
                                stage1_has_we     <= w_stage1_has_we;
                                stage1_has_mem    <= w_stage1_has_mem;
                                stage1_has_mem_we <= w_stage1_has_mem_we;
                                //stage1_alu_op     <= w_stage1_alu_op;
                                stage1_halt       <= w_stage1_halt;

                                d_valid <= f_valid;
                        end else begin
                                d_valid <= 0;
                        end
                        
                                
                        stage1_alu_d  <= w_stage1_alu_d;
                        stage1_alu_d2 <= reg_rd1;
                        e_valid       <= d_valid;
                        valid_stage1  <= d_valid;
                end
                
        end

        // Calculate rd3 data for ALU
        reg [15:0] stage1_rd3;
        always @(*) begin
                stage1_rd3 = 0;
                if (!stall) begin
                        if ((w_stage1_op == `VMICRO16_OP_SW) || (w_stage1_op == `VMICRO16_OP_LW)) begin
                                stage1_rd3 = reg_rd2 + { {11{w_stage1_imm8[4]}}, w_stage1_simm5 };
                                $display($time, "\t\tALU: SWLW: = %d", stage1_rd3);
                        end
                        else if(w_stage1_has_imm8) 
                                stage1_rd3 = { {8{w_stage1_imm8[7]}}, w_stage1_imm8 };
                        else if ((w_stage1_op == `VMICRO16_OP_ARITH_U && stage1_instr[4] == 0)) begin
                                stage1_rd3 = reg_rd2 + { {12{1'b0}}, stage1_instr[3:0] };
                                $display($time, "\t\tALU: ARITH_U: %d + %d = %d", 
                                        reg_rd2, { {12{1'b0}}, stage1_instr[3:0] }, stage1_rd3);
                        end
                        else if ((w_stage1_op == `VMICRO16_OP_ARITH_S && stage1_instr[4] == 0))
                                stage1_rd3 = reg_rd2 + { {12{stage1_instr[3]}}, stage1_instr[3:0] };
                        else
                                stage1_rd3 = reg_rd2;
                end
        end

        wire [4:0]  w_stage1_op;
        wire [7:0]  w_stage1_imm8;
        wire [7:0]  w_stage1_simm5;
        wire        w_stage1_has_imm8;
        wire        w_stage1_has_br;
        wire        w_stage1_has_we;
        wire        w_stage1_has_mem;
        wire        w_stage1_has_mem_we;
        wire [4:0]  w_stage1_alu_op;
        wire [15:0]  w_stage1_alu_d;
        wire        w_stage1_halt;
        vmicro16_dec decoder (
                .instr          (stage1_instr),
                .opcode         (w_stage1_op),
                .rd             (stage1_rs1),
                .ra             (stage1_rs2),
                .imm8           (w_stage1_imm8),
                .simm5          (w_stage1_simm5),
                .has_imm8       (w_stage1_has_imm8   ),
                //.simm5          (w_stage1_simm5      ),
                .has_br         (w_stage1_has_br     ),
                .has_we         (w_stage1_has_we     ),
                //.has_bad       w(stage1_has_bad     ),
                .has_mem        (w_stage1_has_mem    ),
                .has_mem_we     (w_stage1_has_mem_we ),
                .alu_op         (w_stage1_alu_op),
                .halt           (w_stage1_halt)
        );

        // ALU
        wire [15:0] alu_q;
        vmicro16_alu alu (
                .op     (w_stage1_alu_op), 
                .d1     (reg_rd1), 
                .d2     (stage1_rd3), 
                .q      (w_stage1_alu_d)
        );
endmodule

module vmicro16_cpu (
        input clk,
        input reset,
        
        // wishbone peripheral master interface
        //   driven by mmu
        output        wb_mosi_stb_o_regs,    // ...
        output        wb_mosi_cyc_o,
        output        wb_mosi_we_o,
        output [15:0] wb_mosi_addr_o,
        output [15:0] wb_mosi_data_o, // seperate data_o and data_i buses
        input  [15:0] wb_miso_data_i, // seperate data_o and data_i buses
        input         wb_miso_ack_i
);
        wire        valid_stage1;
        wire [4:0]  stage1_op;
        wire [2:0]  stage1_rs1c;
        wire [2:0]  stage1_rs2c;
        wire        stage1_has_imm8;
        wire        stage1_has_br;
        wire        stage1_has_we;
        wire        stage1_has_mem;
        wire        stage1_has_mem_we;
        //wire        stage1_has_bad;
        wire [15:0] stage1_alu_d;
        wire [15:0] stage1_alu_d2;
        wire [15:0] stage1_pc;

        wire [2:0]  reg_rs1;
        wire [2:0]  reg_rs2;
        wire [15:0] reg_rd1;
        wire [15:0] reg_rd2;
        wire [15:0] wb_jmp_target;

        wire        wb_we;
        wire        wb_we_w = reset ? 1'b0 : (wb_we && valid_wb);
        //wire        wb_we_w = 0;
        wire [2:0]  wb_rs1;
        wire [15:0] wb_d;
        vmicro16_regs # (
                .CELL_WIDTH(16),
                .CELL_DEPTH(8)
        ) regs (
                .clk    (clk), 
                .reset  (reset),

                .rs1    (reg_rs1),
                .rd1    (reg_rd1),

                .rs2    (reg_rs2),
                .rd2    (reg_rd2),
                
                .we     (wb_we_w),
                .ws1    (wb_rs1),
                .wd     (wb_d)
        );

        reg jmping = 0;

        wire nop          = !(|stage1_op);
        wire stall_stage1 = (!nop && valid_stage1);
        wire stall_mewb   = (!nop && valid_mewb) && ((stage1_rs1c == mewb_rs1) || ((~stage1_has_imm8) && (stage1_rs2c == mewb_rs1)));
        wire stall_wb     = (!nop && valid_wb)   && ((stage1_rs1c == wb_rs1)   || ((~stage1_has_imm8) && (stage1_rs2c == wb_rs1)));
        //wire stall_mem    = 1'b0;
        wire stall        = |{ stall_stage1,
                               stall_mewb, 
                               stall_wb, 
                               stage1_halt
                               //!mem_valid 
                               };
        
        //reg stall;
        //always @(*) begin
        //        stall = 0;
        //        if (valid_stage1 && |stage1_op)
        //end

        // Stage1
        vmicro16_stage1new stage1 (
                .clk                    (clk), 
                .reset                  (reset), 
                // control signals
                .stall                  (stall), 
                .valid_stage1           (valid_stage1),

                // sync outputs
                .stage1_pc              (stage1_pc), 
                
                // sync decoder outputs
                .stage1_op              (stage1_op), 
                .stage1_rs1c            (stage1_rs1c), 
                .stage1_rs2c            (stage1_rs2c), 
                //.stage1_simm5           (stage1_simm5), 
                .stage1_has_imm8        (stage1_has_imm8),
                .stage1_has_we          (stage1_has_we), 
                .stage1_has_mem         (stage1_has_mem), 
                .stage1_has_br          (stage1_has_br), 
                .stage1_has_mem_we      (stage1_has_mem_we), 
                .stage1_halt            (stage1_halt), 

                // sync alu outputs
                .stage1_alu_d           (stage1_alu_d),
                .stage1_alu_d2          (stage1_alu_d2),

                // Async outputs
                .stage1_rs1             (reg_rs1), 
                .stage1_rs2             (reg_rs2), 
                // Async inputs
                .reg_rd1                (reg_rd1), 
                .reg_rd2                (reg_rd2)
        );

        
        //*
        wire [15:0] mem_out;
        //                     If SW, use calculated address
        wire [15:0] mem_addr = stage1_has_mem ? stage1_alu_d : 16'h00;
        //                     If SW, use register value
        wire [15:0] mem_in   = stage1_has_mem ? stage1_alu_d2 : stage1_alu_d;
        wire        mem_we   = reset ? 1'b0 : (stage1_has_mem_we & valid_stage1);
        wire [1:0]  mem_whl  = 2'b00; // TODO: implement in ISA
        vmicro16_mmu mmu (
                .clk            (clk), 
                .reset          (reset), 

                .req            (stage1_has_mem && valid_stage1),
                .valid          (valid_mem),

                .mem_addr       (mem_addr), 
                .mem_in         (mem_in), 
                .mem_we         (mem_we), 
                .mem_whl        (mem_whl),
                .mem_out        (mem_out),

                // wishbone master interface
                // TODO: Add to top level cpu
                .wb_mosi_stb_o_regs (wb_mosi_stb_o_regs),
                .wb_mosi_cyc_o      (wb_mosi_cyc_o),
                .wb_mosi_we_o       (wb_mosi_we_o),
                .wb_mosi_addr_o     (wb_mosi_addr_o),
                .wb_mosi_data_o     (wb_mosi_data_o),
                .wb_miso_data_i     (wb_miso_data_i),
                .wb_miso_ack_i      (wb_miso_ack_i)
        );

        wire [15:0] mewb_pc;
        wire [15:0] mewb_d;
        wire [15:0] mewb_d2;
        wire [2:0]  mewb_rs1;
        wire [15:0] mewb_jmp_target;
        wire        mewb_has_mem;
        wire        mewb_has_mem_we;
        wire        mewb_has_br;
        wire        mewb_has_we;
        wire        valid_mewb;
        vmicro16_mewb stage_mewb (
                .clk             (clk), 
                .reset           (reset), 

                .valid_stage1    (valid_stage1), 
                .valid_mewb      (valid_mewb),
                .valid_mem       (valid_mem),

                .jmping          (jmping),

                .mem_out         (mem_out), 

                .exme_pc         (stage1_pc), 
                .mewb_pc         (mewb_pc), 

                .exme_d          (stage1_alu_d), 
                .mewb_d          (mewb_d), 
                .exme_d2         (stage1_alu_d2), 
                .mewb_d2         (mewb_d2), 

                .exme_rs1        (stage1_rs1c), 
                .mewb_rs1        (mewb_rs1), 

                .exme_jmp_target (stage1_jmp_target), 
                .mewb_jmp_target (mewb_jmp_target), 

                .exme_has_br     (stage1_has_br), 
                .mewb_has_br     (mewb_has_br), 
                .exme_has_we     (stage1_has_we), 
                .mewb_has_we     (mewb_has_we),  
                .exme_has_mem    (stage1_has_mem), 
                .mewb_has_mem    (mewb_has_mem), 
                .exme_has_mem_we (stage1_has_mem_we), 
                .mewb_has_mem_we (mewb_has_mem_we)
        );

        
        // WB stage
        vmicro16_wb stage_wb (
                .clk             (clk), 
                .reset           (reset), 

                .mewb_d          (mewb_d), 
                .wb_d            (wb_d), 

                .mewb_rs1        (mewb_rs1), 
                .wb_rs1          (wb_rs1), 

                .mewb_has_we     (mewb_has_we), 
                .wb_we           (wb_we), 

                .mewb_has_br     (mewb_has_br), 
                .wb_has_br       (wb_has_br), 

                .mewb_jmp_target (mewb_jmp_target), 
                .wb_jmp_target   (wb_jmp_target), 

                .jmping          (jmping), 

                .valid_mewb      (valid_mewb), 
                .valid_wb        (valid_wb)
        );
endmodule
